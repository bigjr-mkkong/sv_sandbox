
package config_pkg;

endpackage
